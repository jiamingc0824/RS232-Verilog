`timescale 1ns / 1ps

module D4to7Decoder(
    input [3:0] q,
    output [6:0] seg
    );

assign seg = (q == 4'h0)? 7'b0000001:
             (q == 4'h1)? 7'b1001111:
             (q == 4'h2)? 7'b0010010:
             (q == 4'h3)? 7'b0000110:
             (q == 4'h4)? 7'b1001100:
             (q == 4'h5)? 7'b0100100:
             (q == 4'h6)? 7'b0100000:
             (q == 4'h7)? 7'b0001111:
             (q == 4'h8)? 7'b0000000:
             (q == 4'h9)? 7'b0000100:
             (q == 4'hA)? 7'b0001000:
             (q == 4'hB)? 7'b1100000:
             (q == 4'hC)? 7'b0110001:
             (q == 4'hD)? 7'b1000010:
             (q == 4'hE)? 7'b0110000:
             (q == 4'hF)? 7'b0111000:
             7'b1111111;
endmodule
