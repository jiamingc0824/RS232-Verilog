`timescale 1ns / 1ps

module D4to7Decoder(
    );


endmodule
