`timescale 1ns / 1ps

module TopLevel(
    );


endmodule
